        others => x"00000000"
    );

begin

    process (clk)
    begin
        if (clk'event and clk = '1') then
            if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
                report "write collision" severity failure;
            end if;
        
            if (from_zpu.memAWriteEnable = '1') then
                ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
                to_zpu.memARead <= from_zpu.memAWrite;
            else
                to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
            end if;
        end if;
    end process;

    process (clk)
    begin
        if (clk'event and clk = '1') then
            if (from_zpu.memBWriteEnable = '1') then
                ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
                to_zpu.memBRead <= from_zpu.memBWrite;
            else
                to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
            end if;
        end if;
    end process;

end arch;

